TESTE TESTE DE PROGRAMAÇÃO
FUNCIONA PELI AMOR DE DEUSSSS