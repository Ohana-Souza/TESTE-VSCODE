TESTE TESTE DE PROGRAMAÇÃO
FUNCIONA PELI AMOR DE DEUSSSS
sera que agora vai???
LKJKLKLK
klçllklklkl
